module virtual_spi_master(
    input logic clk,
    spi_if.mst_port spi_port
);
    logic [31:0] cnt = '0;
    logic vir_clk = 0;;
    logic [31:0] index_1 = '0;
    logic [3:0] index_2 = 4'hf;

    logic [15:0] mem[0:2000];

    always_ff @(posedge clk) begin
        if(cnt == 32'h0000_0050) begin
            vir_clk <= ~vir_clk;
            cnt <= '0;
        end else begin
            vir_clk <= vir_clk;
            cnt <= cnt + 1;
        end
        mem[0] <= 16'h0555;
        mem[1] <= 16'h1001;
        mem[2] <= 16'h0020;
        mem[3] <= 16'h1002;
        mem[4] <= 16'h0020;
        mem[5] <= 16'h4000;
mem[6] <= 16'h0000;
mem[7] <= 16'h0001;
mem[8] <= 16'h0002;
mem[9] <= 16'h0003;
mem[10] <= 16'h0004;
mem[11] <= 16'h0005;
mem[12] <= 16'h0006;
mem[13] <= 16'h0007;
mem[14] <= 16'h0008;
mem[15] <= 16'h0009;
mem[16] <= 16'h000a;
mem[17] <= 16'h000b;
mem[18] <= 16'h000c;
mem[19] <= 16'h000d;
mem[20] <= 16'h000e;
mem[21] <= 16'h000f;
mem[22] <= 16'h0010;
mem[23] <= 16'h0011;
mem[24] <= 16'h0012;
mem[25] <= 16'h0013;
mem[26] <= 16'h0014;
mem[27] <= 16'h0015;
mem[28] <= 16'h0016;
mem[29] <= 16'h0017;
mem[30] <= 16'h0018;
mem[31] <= 16'h0019;
mem[32] <= 16'h001a;
mem[33] <= 16'h001b;
mem[34] <= 16'h001c;
mem[35] <= 16'h001d;
mem[36] <= 16'h001e;
mem[37] <= 16'h001f;
mem[38] <= 16'h5000;
mem[39] <= 16'h0000;
mem[40] <= 16'h0000;
mem[41] <= 16'h0000;
mem[42] <= 16'h0000;
mem[43] <= 16'h0000;
mem[44] <= 16'h0000;
mem[45] <= 16'h0000;
mem[46] <= 16'h0000;
mem[47] <= 16'h0000;
mem[48] <= 16'h0000;
mem[49] <= 16'h0000;
mem[50] <= 16'h0000;
mem[51] <= 16'h0000;
mem[52] <= 16'h0000;
mem[53] <= 16'h0000;
mem[54] <= 16'h0000;
mem[55] <= 16'h0000;
mem[56] <= 16'h0000;
mem[57] <= 16'h0000;
mem[58] <= 16'h0000;
mem[59] <= 16'h0000;
mem[60] <= 16'h0000;
mem[61] <= 16'h0000;
mem[62] <= 16'h0000;
mem[63] <= 16'h0000;
mem[64] <= 16'h0000;
mem[65] <= 16'h0000;
mem[66] <= 16'h0000;
mem[67] <= 16'h0000;
mem[68] <= 16'h0000;
mem[69] <= 16'h0000;
mem[70] <= 16'h0000;
mem[71] <= 16'h0001;
mem[72] <= 16'h0001;
mem[73] <= 16'h0001;
mem[74] <= 16'h0001;
mem[75] <= 16'h0001;
mem[76] <= 16'h0001;
mem[77] <= 16'h0001;
mem[78] <= 16'h0001;
mem[79] <= 16'h0001;
mem[80] <= 16'h0001;
mem[81] <= 16'h0001;
mem[82] <= 16'h0001;
mem[83] <= 16'h0001;
mem[84] <= 16'h0001;
mem[85] <= 16'h0001;
mem[86] <= 16'h0001;
mem[87] <= 16'h0001;
mem[88] <= 16'h0001;
mem[89] <= 16'h0001;
mem[90] <= 16'h0001;
mem[91] <= 16'h0001;
mem[92] <= 16'h0001;
mem[93] <= 16'h0001;
mem[94] <= 16'h0001;
mem[95] <= 16'h0001;
mem[96] <= 16'h0001;
mem[97] <= 16'h0001;
mem[98] <= 16'h0001;
mem[99] <= 16'h0001;
mem[100] <= 16'h0001;
mem[101] <= 16'h0001;
mem[102] <= 16'h0001;
mem[103] <= 16'h0002;
mem[104] <= 16'h0002;
mem[105] <= 16'h0002;
mem[106] <= 16'h0002;
mem[107] <= 16'h0002;
mem[108] <= 16'h0002;
mem[109] <= 16'h0002;
mem[110] <= 16'h0002;
mem[111] <= 16'h0002;
mem[112] <= 16'h0002;
mem[113] <= 16'h0002;
mem[114] <= 16'h0002;
mem[115] <= 16'h0002;
mem[116] <= 16'h0002;
mem[117] <= 16'h0002;
mem[118] <= 16'h0002;
mem[119] <= 16'h0002;
mem[120] <= 16'h0002;
mem[121] <= 16'h0002;
mem[122] <= 16'h0002;
mem[123] <= 16'h0002;
mem[124] <= 16'h0002;
mem[125] <= 16'h0002;
mem[126] <= 16'h0002;
mem[127] <= 16'h0002;
mem[128] <= 16'h0002;
mem[129] <= 16'h0002;
mem[130] <= 16'h0002;
mem[131] <= 16'h0002;
mem[132] <= 16'h0002;
mem[133] <= 16'h0002;
mem[134] <= 16'h0002;
mem[135] <= 16'h0003;
mem[136] <= 16'h0003;
mem[137] <= 16'h0003;
mem[138] <= 16'h0003;
mem[139] <= 16'h0003;
mem[140] <= 16'h0003;
mem[141] <= 16'h0003;
mem[142] <= 16'h0003;
mem[143] <= 16'h0003;
mem[144] <= 16'h0003;
mem[145] <= 16'h0003;
mem[146] <= 16'h0003;
mem[147] <= 16'h0003;
mem[148] <= 16'h0003;
mem[149] <= 16'h0003;
mem[150] <= 16'h0003;
mem[151] <= 16'h0003;
mem[152] <= 16'h0003;
mem[153] <= 16'h0003;
mem[154] <= 16'h0003;
mem[155] <= 16'h0003;
mem[156] <= 16'h0003;
mem[157] <= 16'h0003;
mem[158] <= 16'h0003;
mem[159] <= 16'h0003;
mem[160] <= 16'h0003;
mem[161] <= 16'h0003;
mem[162] <= 16'h0003;
mem[163] <= 16'h0003;
mem[164] <= 16'h0003;
mem[165] <= 16'h0003;
mem[166] <= 16'h0003;
mem[167] <= 16'h0004;
mem[168] <= 16'h0004;
mem[169] <= 16'h0004;
mem[170] <= 16'h0004;
mem[171] <= 16'h0004;
mem[172] <= 16'h0004;
mem[173] <= 16'h0004;
mem[174] <= 16'h0004;
mem[175] <= 16'h0004;
mem[176] <= 16'h0004;
mem[177] <= 16'h0004;
mem[178] <= 16'h0004;
mem[179] <= 16'h0004;
mem[180] <= 16'h0004;
mem[181] <= 16'h0004;
mem[182] <= 16'h0004;
mem[183] <= 16'h0004;
mem[184] <= 16'h0004;
mem[185] <= 16'h0004;
mem[186] <= 16'h0004;
mem[187] <= 16'h0004;
mem[188] <= 16'h0004;
mem[189] <= 16'h0004;
mem[190] <= 16'h0004;
mem[191] <= 16'h0004;
mem[192] <= 16'h0004;
mem[193] <= 16'h0004;
mem[194] <= 16'h0004;
mem[195] <= 16'h0004;
mem[196] <= 16'h0004;
mem[197] <= 16'h0004;
mem[198] <= 16'h0004;
mem[199] <= 16'h0005;
mem[200] <= 16'h0005;
mem[201] <= 16'h0005;
mem[202] <= 16'h0005;
mem[203] <= 16'h0005;
mem[204] <= 16'h0005;
mem[205] <= 16'h0005;
mem[206] <= 16'h0005;
mem[207] <= 16'h0005;
mem[208] <= 16'h0005;
mem[209] <= 16'h0005;
mem[210] <= 16'h0005;
mem[211] <= 16'h0005;
mem[212] <= 16'h0005;
mem[213] <= 16'h0005;
mem[214] <= 16'h0005;
mem[215] <= 16'h0005;
mem[216] <= 16'h0005;
mem[217] <= 16'h0005;
mem[218] <= 16'h0005;
mem[219] <= 16'h0005;
mem[220] <= 16'h0005;
mem[221] <= 16'h0005;
mem[222] <= 16'h0005;
mem[223] <= 16'h0005;
mem[224] <= 16'h0005;
mem[225] <= 16'h0005;
mem[226] <= 16'h0005;
mem[227] <= 16'h0005;
mem[228] <= 16'h0005;
mem[229] <= 16'h0005;
mem[230] <= 16'h0005;
mem[231] <= 16'h0006;
mem[232] <= 16'h0006;
mem[233] <= 16'h0006;
mem[234] <= 16'h0006;
mem[235] <= 16'h0006;
mem[236] <= 16'h0006;
mem[237] <= 16'h0006;
mem[238] <= 16'h0006;
mem[239] <= 16'h0006;
mem[240] <= 16'h0006;
mem[241] <= 16'h0006;
mem[242] <= 16'h0006;
mem[243] <= 16'h0006;
mem[244] <= 16'h0006;
mem[245] <= 16'h0006;
mem[246] <= 16'h0006;
mem[247] <= 16'h0006;
mem[248] <= 16'h0006;
mem[249] <= 16'h0006;
mem[250] <= 16'h0006;
mem[251] <= 16'h0006;
mem[252] <= 16'h0006;
mem[253] <= 16'h0006;
mem[254] <= 16'h0006;
mem[255] <= 16'h0006;
mem[256] <= 16'h0006;
mem[257] <= 16'h0006;
mem[258] <= 16'h0006;
mem[259] <= 16'h0006;
mem[260] <= 16'h0006;
mem[261] <= 16'h0006;
mem[262] <= 16'h0006;
mem[263] <= 16'h0007;
mem[264] <= 16'h0007;
mem[265] <= 16'h0007;
mem[266] <= 16'h0007;
mem[267] <= 16'h0007;
mem[268] <= 16'h0007;
mem[269] <= 16'h0007;
mem[270] <= 16'h0007;
mem[271] <= 16'h0007;
mem[272] <= 16'h0007;
mem[273] <= 16'h0007;
mem[274] <= 16'h0007;
mem[275] <= 16'h0007;
mem[276] <= 16'h0007;
mem[277] <= 16'h0007;
mem[278] <= 16'h0007;
mem[279] <= 16'h0007;
mem[280] <= 16'h0007;
mem[281] <= 16'h0007;
mem[282] <= 16'h0007;
mem[283] <= 16'h0007;
mem[284] <= 16'h0007;
mem[285] <= 16'h0007;
mem[286] <= 16'h0007;
mem[287] <= 16'h0007;
mem[288] <= 16'h0007;
mem[289] <= 16'h0007;
mem[290] <= 16'h0007;
mem[291] <= 16'h0007;
mem[292] <= 16'h0007;
mem[293] <= 16'h0007;
mem[294] <= 16'h0007;
mem[295] <= 16'h0008;
mem[296] <= 16'h0008;
mem[297] <= 16'h0008;
mem[298] <= 16'h0008;
mem[299] <= 16'h0008;
mem[300] <= 16'h0008;
mem[301] <= 16'h0008;
mem[302] <= 16'h0008;
mem[303] <= 16'h0008;
mem[304] <= 16'h0008;
mem[305] <= 16'h0008;
mem[306] <= 16'h0008;
mem[307] <= 16'h0008;
mem[308] <= 16'h0008;
mem[309] <= 16'h0008;
mem[310] <= 16'h0008;
mem[311] <= 16'h0008;
mem[312] <= 16'h0008;
mem[313] <= 16'h0008;
mem[314] <= 16'h0008;
mem[315] <= 16'h0008;
mem[316] <= 16'h0008;
mem[317] <= 16'h0008;
mem[318] <= 16'h0008;
mem[319] <= 16'h0008;
mem[320] <= 16'h0008;
mem[321] <= 16'h0008;
mem[322] <= 16'h0008;
mem[323] <= 16'h0008;
mem[324] <= 16'h0008;
mem[325] <= 16'h0008;
mem[326] <= 16'h0008;
mem[327] <= 16'h0009;
mem[328] <= 16'h0009;
mem[329] <= 16'h0009;
mem[330] <= 16'h0009;
mem[331] <= 16'h0009;
mem[332] <= 16'h0009;
mem[333] <= 16'h0009;
mem[334] <= 16'h0009;
mem[335] <= 16'h0009;
mem[336] <= 16'h0009;
mem[337] <= 16'h0009;
mem[338] <= 16'h0009;
mem[339] <= 16'h0009;
mem[340] <= 16'h0009;
mem[341] <= 16'h0009;
mem[342] <= 16'h0009;
mem[343] <= 16'h0009;
mem[344] <= 16'h0009;
mem[345] <= 16'h0009;
mem[346] <= 16'h0009;
mem[347] <= 16'h0009;
mem[348] <= 16'h0009;
mem[349] <= 16'h0009;
mem[350] <= 16'h0009;
mem[351] <= 16'h0009;
mem[352] <= 16'h0009;
mem[353] <= 16'h0009;
mem[354] <= 16'h0009;
mem[355] <= 16'h0009;
mem[356] <= 16'h0009;
mem[357] <= 16'h0009;
mem[358] <= 16'h0009;
mem[359] <= 16'h000a;
mem[360] <= 16'h000a;
mem[361] <= 16'h000a;
mem[362] <= 16'h000a;
mem[363] <= 16'h000a;
mem[364] <= 16'h000a;
mem[365] <= 16'h000a;
mem[366] <= 16'h000a;
mem[367] <= 16'h000a;
mem[368] <= 16'h000a;
mem[369] <= 16'h000a;
mem[370] <= 16'h000a;
mem[371] <= 16'h000a;
mem[372] <= 16'h000a;
mem[373] <= 16'h000a;
mem[374] <= 16'h000a;
mem[375] <= 16'h000a;
mem[376] <= 16'h000a;
mem[377] <= 16'h000a;
mem[378] <= 16'h000a;
mem[379] <= 16'h000a;
mem[380] <= 16'h000a;
mem[381] <= 16'h000a;
mem[382] <= 16'h000a;
mem[383] <= 16'h000a;
mem[384] <= 16'h000a;
mem[385] <= 16'h000a;
mem[386] <= 16'h000a;
mem[387] <= 16'h000a;
mem[388] <= 16'h000a;
mem[389] <= 16'h000a;
mem[390] <= 16'h000a;
mem[391] <= 16'h000b;
mem[392] <= 16'h000b;
mem[393] <= 16'h000b;
mem[394] <= 16'h000b;
mem[395] <= 16'h000b;
mem[396] <= 16'h000b;
mem[397] <= 16'h000b;
mem[398] <= 16'h000b;
mem[399] <= 16'h000b;
mem[400] <= 16'h000b;
mem[401] <= 16'h000b;
mem[402] <= 16'h000b;
mem[403] <= 16'h000b;
mem[404] <= 16'h000b;
mem[405] <= 16'h000b;
mem[406] <= 16'h000b;
mem[407] <= 16'h000b;
mem[408] <= 16'h000b;
mem[409] <= 16'h000b;
mem[410] <= 16'h000b;
mem[411] <= 16'h000b;
mem[412] <= 16'h000b;
mem[413] <= 16'h000b;
mem[414] <= 16'h000b;
mem[415] <= 16'h000b;
mem[416] <= 16'h000b;
mem[417] <= 16'h000b;
mem[418] <= 16'h000b;
mem[419] <= 16'h000b;
mem[420] <= 16'h000b;
mem[421] <= 16'h000b;
mem[422] <= 16'h000b;
mem[423] <= 16'h000c;
mem[424] <= 16'h000c;
mem[425] <= 16'h000c;
mem[426] <= 16'h000c;
mem[427] <= 16'h000c;
mem[428] <= 16'h000c;
mem[429] <= 16'h000c;
mem[430] <= 16'h000c;
mem[431] <= 16'h000c;
mem[432] <= 16'h000c;
mem[433] <= 16'h000c;
mem[434] <= 16'h000c;
mem[435] <= 16'h000c;
mem[436] <= 16'h000c;
mem[437] <= 16'h000c;
mem[438] <= 16'h000c;
mem[439] <= 16'h000c;
mem[440] <= 16'h000c;
mem[441] <= 16'h000c;
mem[442] <= 16'h000c;
mem[443] <= 16'h000c;
mem[444] <= 16'h000c;
mem[445] <= 16'h000c;
mem[446] <= 16'h000c;
mem[447] <= 16'h000c;
mem[448] <= 16'h000c;
mem[449] <= 16'h000c;
mem[450] <= 16'h000c;
mem[451] <= 16'h000c;
mem[452] <= 16'h000c;
mem[453] <= 16'h000c;
mem[454] <= 16'h000c;
mem[455] <= 16'h000d;
mem[456] <= 16'h000d;
mem[457] <= 16'h000d;
mem[458] <= 16'h000d;
mem[459] <= 16'h000d;
mem[460] <= 16'h000d;
mem[461] <= 16'h000d;
mem[462] <= 16'h000d;
mem[463] <= 16'h000d;
mem[464] <= 16'h000d;
mem[465] <= 16'h000d;
mem[466] <= 16'h000d;
mem[467] <= 16'h000d;
mem[468] <= 16'h000d;
mem[469] <= 16'h000d;
mem[470] <= 16'h000d;
mem[471] <= 16'h000d;
mem[472] <= 16'h000d;
mem[473] <= 16'h000d;
mem[474] <= 16'h000d;
mem[475] <= 16'h000d;
mem[476] <= 16'h000d;
mem[477] <= 16'h000d;
mem[478] <= 16'h000d;
mem[479] <= 16'h000d;
mem[480] <= 16'h000d;
mem[481] <= 16'h000d;
mem[482] <= 16'h000d;
mem[483] <= 16'h000d;
mem[484] <= 16'h000d;
mem[485] <= 16'h000d;
mem[486] <= 16'h000d;
mem[487] <= 16'h000e;
mem[488] <= 16'h000e;
mem[489] <= 16'h000e;
mem[490] <= 16'h000e;
mem[491] <= 16'h000e;
mem[492] <= 16'h000e;
mem[493] <= 16'h000e;
mem[494] <= 16'h000e;
mem[495] <= 16'h000e;
mem[496] <= 16'h000e;
mem[497] <= 16'h000e;
mem[498] <= 16'h000e;
mem[499] <= 16'h000e;
mem[500] <= 16'h000e;
mem[501] <= 16'h000e;
mem[502] <= 16'h000e;
mem[503] <= 16'h000e;
mem[504] <= 16'h000e;
mem[505] <= 16'h000e;
mem[506] <= 16'h000e;
mem[507] <= 16'h000e;
mem[508] <= 16'h000e;
mem[509] <= 16'h000e;
mem[510] <= 16'h000e;
mem[511] <= 16'h000e;
mem[512] <= 16'h000e;
mem[513] <= 16'h000e;
mem[514] <= 16'h000e;
mem[515] <= 16'h000e;
mem[516] <= 16'h000e;
mem[517] <= 16'h000e;
mem[518] <= 16'h000e;
mem[519] <= 16'h000f;
mem[520] <= 16'h000f;
mem[521] <= 16'h000f;
mem[522] <= 16'h000f;
mem[523] <= 16'h000f;
mem[524] <= 16'h000f;
mem[525] <= 16'h000f;
mem[526] <= 16'h000f;
mem[527] <= 16'h000f;
mem[528] <= 16'h000f;
mem[529] <= 16'h000f;
mem[530] <= 16'h000f;
mem[531] <= 16'h000f;
mem[532] <= 16'h000f;
mem[533] <= 16'h000f;
mem[534] <= 16'h000f;
mem[535] <= 16'h000f;
mem[536] <= 16'h000f;
mem[537] <= 16'h000f;
mem[538] <= 16'h000f;
mem[539] <= 16'h000f;
mem[540] <= 16'h000f;
mem[541] <= 16'h000f;
mem[542] <= 16'h000f;
mem[543] <= 16'h000f;
mem[544] <= 16'h000f;
mem[545] <= 16'h000f;
mem[546] <= 16'h000f;
mem[547] <= 16'h000f;
mem[548] <= 16'h000f;
mem[549] <= 16'h000f;
mem[550] <= 16'h000f;
mem[551] <= 16'h0010;
mem[552] <= 16'h0010;
mem[553] <= 16'h0010;
mem[554] <= 16'h0010;
mem[555] <= 16'h0010;
mem[556] <= 16'h0010;
mem[557] <= 16'h0010;
mem[558] <= 16'h0010;
mem[559] <= 16'h0010;
mem[560] <= 16'h0010;
mem[561] <= 16'h0010;
mem[562] <= 16'h0010;
mem[563] <= 16'h0010;
mem[564] <= 16'h0010;
mem[565] <= 16'h0010;
mem[566] <= 16'h0010;
mem[567] <= 16'h0010;
mem[568] <= 16'h0010;
mem[569] <= 16'h0010;
mem[570] <= 16'h0010;
mem[571] <= 16'h0010;
mem[572] <= 16'h0010;
mem[573] <= 16'h0010;
mem[574] <= 16'h0010;
mem[575] <= 16'h0010;
mem[576] <= 16'h0010;
mem[577] <= 16'h0010;
mem[578] <= 16'h0010;
mem[579] <= 16'h0010;
mem[580] <= 16'h0010;
mem[581] <= 16'h0010;
mem[582] <= 16'h0010;
mem[583] <= 16'h0011;
mem[584] <= 16'h0011;
mem[585] <= 16'h0011;
mem[586] <= 16'h0011;
mem[587] <= 16'h0011;
mem[588] <= 16'h0011;
mem[589] <= 16'h0011;
mem[590] <= 16'h0011;
mem[591] <= 16'h0011;
mem[592] <= 16'h0011;
mem[593] <= 16'h0011;
mem[594] <= 16'h0011;
mem[595] <= 16'h0011;
mem[596] <= 16'h0011;
mem[597] <= 16'h0011;
mem[598] <= 16'h0011;
mem[599] <= 16'h0011;
mem[600] <= 16'h0011;
mem[601] <= 16'h0011;
mem[602] <= 16'h0011;
mem[603] <= 16'h0011;
mem[604] <= 16'h0011;
mem[605] <= 16'h0011;
mem[606] <= 16'h0011;
mem[607] <= 16'h0011;
mem[608] <= 16'h0011;
mem[609] <= 16'h0011;
mem[610] <= 16'h0011;
mem[611] <= 16'h0011;
mem[612] <= 16'h0011;
mem[613] <= 16'h0011;
mem[614] <= 16'h0011;
mem[615] <= 16'h0012;
mem[616] <= 16'h0012;
mem[617] <= 16'h0012;
mem[618] <= 16'h0012;
mem[619] <= 16'h0012;
mem[620] <= 16'h0012;
mem[621] <= 16'h0012;
mem[622] <= 16'h0012;
mem[623] <= 16'h0012;
mem[624] <= 16'h0012;
mem[625] <= 16'h0012;
mem[626] <= 16'h0012;
mem[627] <= 16'h0012;
mem[628] <= 16'h0012;
mem[629] <= 16'h0012;
mem[630] <= 16'h0012;
mem[631] <= 16'h0012;
mem[632] <= 16'h0012;
mem[633] <= 16'h0012;
mem[634] <= 16'h0012;
mem[635] <= 16'h0012;
mem[636] <= 16'h0012;
mem[637] <= 16'h0012;
mem[638] <= 16'h0012;
mem[639] <= 16'h0012;
mem[640] <= 16'h0012;
mem[641] <= 16'h0012;
mem[642] <= 16'h0012;
mem[643] <= 16'h0012;
mem[644] <= 16'h0012;
mem[645] <= 16'h0012;
mem[646] <= 16'h0012;
mem[647] <= 16'h0013;
mem[648] <= 16'h0013;
mem[649] <= 16'h0013;
mem[650] <= 16'h0013;
mem[651] <= 16'h0013;
mem[652] <= 16'h0013;
mem[653] <= 16'h0013;
mem[654] <= 16'h0013;
mem[655] <= 16'h0013;
mem[656] <= 16'h0013;
mem[657] <= 16'h0013;
mem[658] <= 16'h0013;
mem[659] <= 16'h0013;
mem[660] <= 16'h0013;
mem[661] <= 16'h0013;
mem[662] <= 16'h0013;
mem[663] <= 16'h0013;
mem[664] <= 16'h0013;
mem[665] <= 16'h0013;
mem[666] <= 16'h0013;
mem[667] <= 16'h0013;
mem[668] <= 16'h0013;
mem[669] <= 16'h0013;
mem[670] <= 16'h0013;
mem[671] <= 16'h0013;
mem[672] <= 16'h0013;
mem[673] <= 16'h0013;
mem[674] <= 16'h0013;
mem[675] <= 16'h0013;
mem[676] <= 16'h0013;
mem[677] <= 16'h0013;
mem[678] <= 16'h0013;
mem[679] <= 16'h0014;
mem[680] <= 16'h0014;
mem[681] <= 16'h0014;
mem[682] <= 16'h0014;
mem[683] <= 16'h0014;
mem[684] <= 16'h0014;
mem[685] <= 16'h0014;
mem[686] <= 16'h0014;
mem[687] <= 16'h0014;
mem[688] <= 16'h0014;
mem[689] <= 16'h0014;
mem[690] <= 16'h0014;
mem[691] <= 16'h0014;
mem[692] <= 16'h0014;
mem[693] <= 16'h0014;
mem[694] <= 16'h0014;
mem[695] <= 16'h0014;
mem[696] <= 16'h0014;
mem[697] <= 16'h0014;
mem[698] <= 16'h0014;
mem[699] <= 16'h0014;
mem[700] <= 16'h0014;
mem[701] <= 16'h0014;
mem[702] <= 16'h0014;
mem[703] <= 16'h0014;
mem[704] <= 16'h0014;
mem[705] <= 16'h0014;
mem[706] <= 16'h0014;
mem[707] <= 16'h0014;
mem[708] <= 16'h0014;
mem[709] <= 16'h0014;
mem[710] <= 16'h0014;
mem[711] <= 16'h0015;
mem[712] <= 16'h0015;
mem[713] <= 16'h0015;
mem[714] <= 16'h0015;
mem[715] <= 16'h0015;
mem[716] <= 16'h0015;
mem[717] <= 16'h0015;
mem[718] <= 16'h0015;
mem[719] <= 16'h0015;
mem[720] <= 16'h0015;
mem[721] <= 16'h0015;
mem[722] <= 16'h0015;
mem[723] <= 16'h0015;
mem[724] <= 16'h0015;
mem[725] <= 16'h0015;
mem[726] <= 16'h0015;
mem[727] <= 16'h0015;
mem[728] <= 16'h0015;
mem[729] <= 16'h0015;
mem[730] <= 16'h0015;
mem[731] <= 16'h0015;
mem[732] <= 16'h0015;
mem[733] <= 16'h0015;
mem[734] <= 16'h0015;
mem[735] <= 16'h0015;
mem[736] <= 16'h0015;
mem[737] <= 16'h0015;
mem[738] <= 16'h0015;
mem[739] <= 16'h0015;
mem[740] <= 16'h0015;
mem[741] <= 16'h0015;
mem[742] <= 16'h0015;
mem[743] <= 16'h0016;
mem[744] <= 16'h0016;
mem[745] <= 16'h0016;
mem[746] <= 16'h0016;
mem[747] <= 16'h0016;
mem[748] <= 16'h0016;
mem[749] <= 16'h0016;
mem[750] <= 16'h0016;
mem[751] <= 16'h0016;
mem[752] <= 16'h0016;
mem[753] <= 16'h0016;
mem[754] <= 16'h0016;
mem[755] <= 16'h0016;
mem[756] <= 16'h0016;
mem[757] <= 16'h0016;
mem[758] <= 16'h0016;
mem[759] <= 16'h0016;
mem[760] <= 16'h0016;
mem[761] <= 16'h0016;
mem[762] <= 16'h0016;
mem[763] <= 16'h0016;
mem[764] <= 16'h0016;
mem[765] <= 16'h0016;
mem[766] <= 16'h0016;
mem[767] <= 16'h0016;
mem[768] <= 16'h0016;
mem[769] <= 16'h0016;
mem[770] <= 16'h0016;
mem[771] <= 16'h0016;
mem[772] <= 16'h0016;
mem[773] <= 16'h0016;
mem[774] <= 16'h0016;
mem[775] <= 16'h0017;
mem[776] <= 16'h0017;
mem[777] <= 16'h0017;
mem[778] <= 16'h0017;
mem[779] <= 16'h0017;
mem[780] <= 16'h0017;
mem[781] <= 16'h0017;
mem[782] <= 16'h0017;
mem[783] <= 16'h0017;
mem[784] <= 16'h0017;
mem[785] <= 16'h0017;
mem[786] <= 16'h0017;
mem[787] <= 16'h0017;
mem[788] <= 16'h0017;
mem[789] <= 16'h0017;
mem[790] <= 16'h0017;
mem[791] <= 16'h0017;
mem[792] <= 16'h0017;
mem[793] <= 16'h0017;
mem[794] <= 16'h0017;
mem[795] <= 16'h0017;
mem[796] <= 16'h0017;
mem[797] <= 16'h0017;
mem[798] <= 16'h0017;
mem[799] <= 16'h0017;
mem[800] <= 16'h0017;
mem[801] <= 16'h0017;
mem[802] <= 16'h0017;
mem[803] <= 16'h0017;
mem[804] <= 16'h0017;
mem[805] <= 16'h0017;
mem[806] <= 16'h0017;
mem[807] <= 16'h0018;
mem[808] <= 16'h0018;
mem[809] <= 16'h0018;
mem[810] <= 16'h0018;
mem[811] <= 16'h0018;
mem[812] <= 16'h0018;
mem[813] <= 16'h0018;
mem[814] <= 16'h0018;
mem[815] <= 16'h0018;
mem[816] <= 16'h0018;
mem[817] <= 16'h0018;
mem[818] <= 16'h0018;
mem[819] <= 16'h0018;
mem[820] <= 16'h0018;
mem[821] <= 16'h0018;
mem[822] <= 16'h0018;
mem[823] <= 16'h0018;
mem[824] <= 16'h0018;
mem[825] <= 16'h0018;
mem[826] <= 16'h0018;
mem[827] <= 16'h0018;
mem[828] <= 16'h0018;
mem[829] <= 16'h0018;
mem[830] <= 16'h0018;
mem[831] <= 16'h0018;
mem[832] <= 16'h0018;
mem[833] <= 16'h0018;
mem[834] <= 16'h0018;
mem[835] <= 16'h0018;
mem[836] <= 16'h0018;
mem[837] <= 16'h0018;
mem[838] <= 16'h0018;
mem[839] <= 16'h0019;
mem[840] <= 16'h0019;
mem[841] <= 16'h0019;
mem[842] <= 16'h0019;
mem[843] <= 16'h0019;
mem[844] <= 16'h0019;
mem[845] <= 16'h0019;
mem[846] <= 16'h0019;
mem[847] <= 16'h0019;
mem[848] <= 16'h0019;
mem[849] <= 16'h0019;
mem[850] <= 16'h0019;
mem[851] <= 16'h0019;
mem[852] <= 16'h0019;
mem[853] <= 16'h0019;
mem[854] <= 16'h0019;
mem[855] <= 16'h0019;
mem[856] <= 16'h0019;
mem[857] <= 16'h0019;
mem[858] <= 16'h0019;
mem[859] <= 16'h0019;
mem[860] <= 16'h0019;
mem[861] <= 16'h0019;
mem[862] <= 16'h0019;
mem[863] <= 16'h0019;
mem[864] <= 16'h0019;
mem[865] <= 16'h0019;
mem[866] <= 16'h0019;
mem[867] <= 16'h0019;
mem[868] <= 16'h0019;
mem[869] <= 16'h0019;
mem[870] <= 16'h0019;
mem[871] <= 16'h001a;
mem[872] <= 16'h001a;
mem[873] <= 16'h001a;
mem[874] <= 16'h001a;
mem[875] <= 16'h001a;
mem[876] <= 16'h001a;
mem[877] <= 16'h001a;
mem[878] <= 16'h001a;
mem[879] <= 16'h001a;
mem[880] <= 16'h001a;
mem[881] <= 16'h001a;
mem[882] <= 16'h001a;
mem[883] <= 16'h001a;
mem[884] <= 16'h001a;
mem[885] <= 16'h001a;
mem[886] <= 16'h001a;
mem[887] <= 16'h001a;
mem[888] <= 16'h001a;
mem[889] <= 16'h001a;
mem[890] <= 16'h001a;
mem[891] <= 16'h001a;
mem[892] <= 16'h001a;
mem[893] <= 16'h001a;
mem[894] <= 16'h001a;
mem[895] <= 16'h001a;
mem[896] <= 16'h001a;
mem[897] <= 16'h001a;
mem[898] <= 16'h001a;
mem[899] <= 16'h001a;
mem[900] <= 16'h001a;
mem[901] <= 16'h001a;
mem[902] <= 16'h001a;
mem[903] <= 16'h001b;
mem[904] <= 16'h001b;
mem[905] <= 16'h001b;
mem[906] <= 16'h001b;
mem[907] <= 16'h001b;
mem[908] <= 16'h001b;
mem[909] <= 16'h001b;
mem[910] <= 16'h001b;
mem[911] <= 16'h001b;
mem[912] <= 16'h001b;
mem[913] <= 16'h001b;
mem[914] <= 16'h001b;
mem[915] <= 16'h001b;
mem[916] <= 16'h001b;
mem[917] <= 16'h001b;
mem[918] <= 16'h001b;
mem[919] <= 16'h001b;
mem[920] <= 16'h001b;
mem[921] <= 16'h001b;
mem[922] <= 16'h001b;
mem[923] <= 16'h001b;
mem[924] <= 16'h001b;
mem[925] <= 16'h001b;
mem[926] <= 16'h001b;
mem[927] <= 16'h001b;
mem[928] <= 16'h001b;
mem[929] <= 16'h001b;
mem[930] <= 16'h001b;
mem[931] <= 16'h001b;
mem[932] <= 16'h001b;
mem[933] <= 16'h001b;
mem[934] <= 16'h001b;
mem[935] <= 16'h001c;
mem[936] <= 16'h001c;
mem[937] <= 16'h001c;
mem[938] <= 16'h001c;
mem[939] <= 16'h001c;
mem[940] <= 16'h001c;
mem[941] <= 16'h001c;
mem[942] <= 16'h001c;
mem[943] <= 16'h001c;
mem[944] <= 16'h001c;
mem[945] <= 16'h001c;
mem[946] <= 16'h001c;
mem[947] <= 16'h001c;
mem[948] <= 16'h001c;
mem[949] <= 16'h001c;
mem[950] <= 16'h001c;
mem[951] <= 16'h001c;
mem[952] <= 16'h001c;
mem[953] <= 16'h001c;
mem[954] <= 16'h001c;
mem[955] <= 16'h001c;
mem[956] <= 16'h001c;
mem[957] <= 16'h001c;
mem[958] <= 16'h001c;
mem[959] <= 16'h001c;
mem[960] <= 16'h001c;
mem[961] <= 16'h001c;
mem[962] <= 16'h001c;
mem[963] <= 16'h001c;
mem[964] <= 16'h001c;
mem[965] <= 16'h001c;
mem[966] <= 16'h001c;
mem[967] <= 16'h001d;
mem[968] <= 16'h001d;
mem[969] <= 16'h001d;
mem[970] <= 16'h001d;
mem[971] <= 16'h001d;
mem[972] <= 16'h001d;
mem[973] <= 16'h001d;
mem[974] <= 16'h001d;
mem[975] <= 16'h001d;
mem[976] <= 16'h001d;
mem[977] <= 16'h001d;
mem[978] <= 16'h001d;
mem[979] <= 16'h001d;
mem[980] <= 16'h001d;
mem[981] <= 16'h001d;
mem[982] <= 16'h001d;
mem[983] <= 16'h001d;
mem[984] <= 16'h001d;
mem[985] <= 16'h001d;
mem[986] <= 16'h001d;
mem[987] <= 16'h001d;
mem[988] <= 16'h001d;
mem[989] <= 16'h001d;
mem[990] <= 16'h001d;
mem[991] <= 16'h001d;
mem[992] <= 16'h001d;
mem[993] <= 16'h001d;
mem[994] <= 16'h001d;
mem[995] <= 16'h001d;
mem[996] <= 16'h001d;
mem[997] <= 16'h001d;
mem[998] <= 16'h001d;
mem[999] <= 16'h001e;
mem[1000] <= 16'h001e;
mem[1001] <= 16'h001e;
mem[1002] <= 16'h001e;
mem[1003] <= 16'h001e;
mem[1004] <= 16'h001e;
mem[1005] <= 16'h001e;
mem[1006] <= 16'h001e;
mem[1007] <= 16'h001e;
mem[1008] <= 16'h001e;
mem[1009] <= 16'h001e;
mem[1010] <= 16'h001e;
mem[1011] <= 16'h001e;
mem[1012] <= 16'h001e;
mem[1013] <= 16'h001e;
mem[1014] <= 16'h001e;
mem[1015] <= 16'h001e;
mem[1016] <= 16'h001e;
mem[1017] <= 16'h001e;
mem[1018] <= 16'h001e;
mem[1019] <= 16'h001e;
mem[1020] <= 16'h001e;
mem[1021] <= 16'h001e;
mem[1022] <= 16'h001e;
mem[1023] <= 16'h001e;
mem[1024] <= 16'h001e;
mem[1025] <= 16'h001e;
mem[1026] <= 16'h001e;
mem[1027] <= 16'h001e;
mem[1028] <= 16'h001e;
mem[1029] <= 16'h001e;
mem[1030] <= 16'h001e;
mem[1031] <= 16'h001f;
mem[1032] <= 16'h001f;
mem[1033] <= 16'h001f;
mem[1034] <= 16'h001f;
mem[1035] <= 16'h001f;
mem[1036] <= 16'h001f;
mem[1037] <= 16'h001f;
mem[1038] <= 16'h001f;
mem[1039] <= 16'h001f;
mem[1040] <= 16'h001f;
mem[1041] <= 16'h001f;
mem[1042] <= 16'h001f;
mem[1043] <= 16'h001f;
mem[1044] <= 16'h001f;
mem[1045] <= 16'h001f;
mem[1046] <= 16'h001f;
mem[1047] <= 16'h001f;
mem[1048] <= 16'h001f;
mem[1049] <= 16'h001f;
mem[1050] <= 16'h001f;
mem[1051] <= 16'h001f;
mem[1052] <= 16'h001f;
mem[1053] <= 16'h001f;
mem[1054] <= 16'h001f;
mem[1055] <= 16'h001f;
mem[1056] <= 16'h001f;
mem[1057] <= 16'h001f;
mem[1058] <= 16'h001f;
mem[1059] <= 16'h001f;
mem[1060] <= 16'h001f;
mem[1061] <= 16'h001f;
mem[1062] <= 16'h001f;
mem[1063] <= 16'h3000;
mem[1064] <= 16'h6000;
mem[1065] <= 16'h0000;
mem[1066] <= 16'h0000;
mem[1067] <= 16'h0000;
mem[1068] <= 16'h0000;
mem[1069] <= 16'h0000;
mem[1070] <= 16'h0000;
mem[1071] <= 16'h0000;
mem[1072] <= 16'h0000;
mem[1073] <= 16'h0000;
mem[1074] <= 16'h0000;
mem[1075] <= 16'h0000;
mem[1076] <= 16'h0000;
mem[1077] <= 16'h0000;
mem[1078] <= 16'h0000;
mem[1079] <= 16'h0000;
mem[1080] <= 16'h0000;
mem[1081] <= 16'h0000;
mem[1082] <= 16'h0000;
mem[1083] <= 16'h0000;
mem[1084] <= 16'h0000;
mem[1085] <= 16'h0000;
mem[1086] <= 16'h0000;
mem[1087] <= 16'h0000;
mem[1088] <= 16'h0000;
mem[1089] <= 16'h0000;
mem[1090] <= 16'h0000;
mem[1091] <= 16'h0000;
mem[1092] <= 16'h0000;
mem[1093] <= 16'h0000;
mem[1094] <= 16'h0000;
mem[1095] <= 16'h0000;
mem[1096] <= 16'h0000;
mem[1097] <= 16'h0000;

    end

    always_ff @(posedge vir_clk) begin
        spi_port.sclk <= ~spi_port.sclk;
    end

    always_ff @(negedge spi_port.sclk) begin
        if(index_2 == 4'h0) begin
            index_2 <= 4'hf;
            index_1 <= index_1 + 1;
        end else begin
            index_2 <= index_2 - 4'h1;
        end
    end
    assign spi_port.mosi = mem[index_1][index_2];


endmodule
