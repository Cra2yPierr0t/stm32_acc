module Controller #(
    parameter ADDR_SIZE = 10,
    parameter WORD_SIZE = 16,
    parameter PE_NUMBER = 64,
    parameter MEM_HEAD_ADDR = 16'h000f,
    parameter ZERO_POINT_ADDR = 16'hffff,
    parameter START_CAL = 4'h3,
    parameter WRITE_VEC = 4'h4,
    parameter WRITE_MAT = 4'h5,
    parameter READ_RESULT = 4'h6
)(
    input   clk,
    bus_if.slv_port spi_2_bus_if,
    output  logic read,
    output  logic reset,
    bus_if.slv_port vec_csr_if,
    bus_if.slv_port mat_csr_if,
    bus_if.slv_port csr_if,
    output  logic [ADDR_SIZE-1:0] pe_t_o_addr[0:PE_NUMBER-1],
    output  logic [ADDR_SIZE-1:0] l_d_o_addr,
    output  logic [WORD_SIZE-1:0] w_data,
    output  logic [ADDR_SIZE-1:0] w_addr,
    output  logic w_en
);

parameter WAIT  = 2'b00;
parameter CAL   = 2'b01;
parameter READ  = 2'b10;

parameter MEM_WAIT  = 2'b00;
parameter MEM_FETCH = 2'b01;
parameter MEM_WRITE = 2'b10;
parameter MEM_CAL_WAIT = 2'b11;

    logic [7:0] row_size;
    logic [7:0] column_size;

    logic [7:0] mem_index = '0;

    logic [7:0] cal_cnt = 8'h00;
    logic [7:0] read_cnt = 8'h00;

    logic [7:0] row_cnt = '0;
    logic [7:0] column_cnt = '0;

    logic   run_req = 0;

    logic [1:0] array_state = WAIT;
    logic [1:0] mem_state   = WAIT;

    logic [ADDR_SIZE-1:0] w_addr_buf = '0;
    logic [ADDR_SIZE-1:0] w_addr_cnt = '0;

    always_ff @(posedge vec_csr_if.valid) begin
        row_size    <= vec_csr_if.data;
    end
    always_ff @(posedge mat_csr_if.valid) begin
        column_size <= mat_csr_if.data;
    end
    always_ff @(posedge csr_if.valid) begin
        run_req <= csr_if.data[0];
    end

    always_ff @(posedge clk) begin
        case(array_state)
            WAIT    : begin
                if(run_req == 1) begin
                    array_state <= CAL;
                end else begin
                    array_state <= WAIT;
                end
                reset   <= 1;
                read    <= 0;
                vec_csr_if.ready <= 1;
                mat_csr_if.ready <= 1;
                csr_if.ready <= 1;
            end
            CAL     : begin
                if(cal_cnt < row_size + column_size - 1) begin
                    cal_cnt <= cal_cnt + 8'h01;
                end else begin
                    array_state   <= READ;
                    cal_cnt <= 8'h00;
                end
                reset   <= 0;
                read    <= 0;
                vec_csr_if.ready <= 0;
                mat_csr_if.ready <= 0;
                csr_if.ready <= 0;
            end
            READ    : begin
                if(read_cnt < column_size - 1) begin //case文でステートマシンを作るときのカスみたいな記述
                    read_cnt <= read_cnt + 8'h01;
                end else begin
                    array_state   <= WAIT;
                    read_cnt <= 8'h00;
                end
                reset   <= 0;
                read    <= 1;
                vec_csr_if.ready <= 0;
                mat_csr_if.ready <= 0;
                csr_if.ready <= 0;
            end
        endcase

        case(mem_state)
            MEM_WAIT    : begin
                if(run_req == 1) begin
                    mem_state <= MEM_FETCH;
                end else begin
                    mem_state <= MEM_WAIT;
                end
                l_d_o_addr <= ZERO_POINT_ADDR;
                //w_en        <= '0;
                w_addr_cnt  <= '0;
            end
            MEM_FETCH   : begin
                if(column_cnt < column_size) begin
                    column_cnt <= column_cnt + 1;
                    mem_index <= mem_index + column_size;
                end else begin
                    column_cnt <= '0;
                    mem_index <= '0;
                end
                if(row_cnt < row_size) begin    //vec fetch
                    l_d_o_addr <= MEM_HEAD_ADDR + row_cnt;
                    row_cnt <= row_cnt + 1;
                    mem_state <= mem_state;
                end else begin
                    l_d_o_addr <= ZERO_POINT_ADDR;
                    row_cnt <= '0;
                    mem_state <= MEM_CAL_WAIT;
                end
            end
            MEM_CAL_WAIT    : begin
                if(cal_cnt < row_size + column_size - 1) begin
                    mem_state <= mem_state;
                end else begin
                    mem_state <= MEM_WRITE;
                end
            end
            MEM_WRITE   : begin
                if(read_cnt < column_size - 1) begin
                    mem_state <= mem_state;
                end else begin
                    mem_state <= MEM_WAIT;
                end
                //w_en        <= '1;
                w_addr      <= w_addr_buf + 1 + w_addr_cnt;
                w_addr_cnt  <= w_addr_cnt + 1;
            end
        endcase
    end
    genvar i;
    generate 
    for(i = 0; i < PE_NUMBER; i = i + 1) begin : gen_fetch_system
        always_ff @(posedge clk) begin
            if(mem_state == MEM_FETCH) begin
                if(row_size > i) begin
                    if(column_cnt < column_size) begin
                        pe_t_o_addr[i]  <= MEM_HEAD_ADDR + row_size + i + mem_index;
                        w_addr_buf      <= MEM_HEAD_ADDR + row_size + i + mem_index;
                    end else begin
                        pe_t_o_addr[i]  <= ZERO_POINT_ADDR;
                        w_addr_buf      <= w_addr_buf;
                    end
                end else begin
                    pe_t_o_addr[i] <= ZERO_POINT_ADDR; 
                end
            end else begin
                pe_t_o_addr[i] <= ZERO_POINT_ADDR; 
            end
        end
    end
    endgenerate

    logic [1:0] spi_shift_reg;
    logic [1:0] vec_shift_reg;
    logic [1:0] mat_shift_reg;

    logic write_vec_flag = 0;
    logic write_mat_flag = 0;

    logic end_vec_flag = 0;
    logic end_mat_flag = 0;

    logic [9:0] mat_sub_cnt = '0;
    logic [9:0] mat_sub_sub_cnt = '0;

    logic [9:0] vec_addr = '0;
    logic [9:0] mat_addr = '0;

    always_ff @(posedge clk) begin
        spi_shift_reg <= {spi_shift_reg[0], spi_2_bus_if.valid};
        vec_shift_reg <= {vec_shift_reg[0], end_vec_flag};
        mat_shift_reg <= {mat_shift_reg[0], end_mat_flag};
        if((write_vec_flag == 0) && (write_mat_flag == 0)) begin
            if(spi_shift_reg == 2'b01) begin
                case(spi_2_bus_if.data[15:12])
                    START_CAL   : begin
                    end
                    WRITE_VEC   : begin
                        write_vec_flag <= 1;
                    end
                    WRITE_MAT   : begin
                        write_mat_flag <= 1;
                    end
                    READ_RESULT : begin
                    end
                    default     : begin
                    end
                endcase
            end else begin
                if(vec_shift_reg == 2'b01) begin
                    write_vec_flag <= 0;
                end
                if(mat_shift_reg == 2'b01) begin
                    write_mat_flag <= 0;
                end
            end
        end

        if(write_vec_flag == 1) begin
            if(spi_shift_reg == 2'b01) begin
                w_en <= 1;
                w_addr <= vec_addr;
                w_data <= spi_2_bus_if.data;
                if(vec_addr == vec_csr_if.data - 1) begin
                    vec_addr <= 0;
                    write_vec_flag <= 0;
                    end_vec_flag <= 1;
                end else begin
                    vec_addr <= vec_addr + 1;
                    end_vec_flag <= 0;
                end
            end else begin
                w_en <= 0;
            end
        end else if(write_mat_flag == 1) begin
            if(spi_shift_reg == 2'b01) begin
                w_en <= 1;
                w_addr <= mat_addr + vec_csr_if.data;
                w_data <= spi_2_bus_if.data;
                if((mat_sub_cnt == mat_csr_if.data - 1) && (mat_sub_sub_cnt == vec_csr_if.data - 1)) begin
                    mat_sub_cnt <= 0;
                    end_mat_flag <= 1;
                    mat_addr <= 0;
                end else if(mat_sub_sub_cnt == vec_csr_if.data - 1) begin
                    mat_sub_sub_cnt <= 0;
                    mat_sub_cnt <= mat_sub_cnt + 1;
                end else begin
                    mat_sub_sub_cnt <= mat_sub_sub_cnt + 1;
                    mat_sub_cnt <= mat_sub_cnt;
                    mat_addr <= mat_addr + 1;
                    end_mat_flag <= 0;
                end
            end else begin
                w_en <= 0;
            end
        end else begin
            w_en <= 0;
            mat_addr <= 0;
            vec_addr <= 0;
        end
    end

endmodule
